library IEEE;
use IEEE.std_logic_1164.all;

-- 16-bit Bus
signal bus : std_logic_vector (15 downto 0);
